package int_types;
   typedef logic [3:0] INT04_t;
   typedef logic [40:0] INT41_t;
endpackage
